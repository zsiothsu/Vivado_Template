`define ADD_NUM 1